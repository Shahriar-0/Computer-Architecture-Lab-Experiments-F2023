module InstructionFetch()