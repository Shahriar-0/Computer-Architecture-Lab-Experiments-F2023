
module WB_Stage(clk, rst);

    parameter N = 32;
    input wire[0:0] clk, rst;

endmodule